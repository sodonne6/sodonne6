module invert1(
input wire d,
output wire notd
    );
    
    assign notd= ~d; //invert bit
endmodule
